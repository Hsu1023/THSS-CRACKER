library verilog;
use verilog.vl_types.all;
entity eda2_vlg_vec_tst is
end eda2_vlg_vec_tst;
