library verilog;
use verilog.vl_types.all;
entity eda1_vlg_vec_tst is
end eda1_vlg_vec_tst;
